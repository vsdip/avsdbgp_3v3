* SPICE3 file created from bgr1.ext - technology: scmos

.option scale=0.1u

M1000 N001 N002 N002 N001 pfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240
M1001 0 N003 N004 0 nfet w=200 l=50
+  ad=6000 pd=1300 as=3909.43 ps=460.377
M1002 N003 N003 N006 0 nfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240
M1003 N005 N003 N002 0 nfet w=100 l=50
+  ad=1892.86 pd=253.571 as=1916.67 ps=258.333
M1004 N002 N004 0 0 nfet w=20 l=20
+  ad=383.333 pd=51.6667 as=600 ps=130
R0 N005 N007 nwellResistor w=12 l=103
M1005 N001 N002 vref N001 pfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240
R1 N001 N004 nwellResistor w=12 l=15428
R2 vref vctat nwellResistor w=12 l=1275
M1006 N003 N002 N001 N001 pfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240
C0 N001 N002 7.36fF
C1 N004 0 2.57fF
C2 N003 0 8.80fF
C3 N001 0 58.37fF
