magic
tech scmos
timestamp 1593517187
<< nwell >>
rect -140 -10 -10 130
rect 10 -10 140 130
rect 160 -10 290 130
<< ntransistor >>
rect -290 -210 -240 -10
rect -190 -50 -170 -30
rect -100 -160 -50 -60
rect 50 -160 100 -60
<< ptransistor >>
rect -100 10 -50 110
rect 50 10 100 110
rect 200 10 250 110
<< ndiffusion >>
rect -310 -15 -290 -10
rect -310 -25 -305 -15
rect -294 -25 -290 -15
rect -310 -35 -290 -25
rect -310 -45 -305 -35
rect -294 -45 -290 -35
rect -310 -55 -290 -45
rect -310 -65 -305 -55
rect -294 -65 -290 -55
rect -310 -75 -290 -65
rect -310 -85 -305 -75
rect -294 -85 -290 -75
rect -310 -95 -290 -85
rect -310 -105 -305 -95
rect -294 -105 -290 -95
rect -310 -115 -290 -105
rect -310 -125 -305 -115
rect -294 -125 -290 -115
rect -310 -135 -290 -125
rect -310 -145 -305 -135
rect -294 -145 -290 -135
rect -310 -155 -290 -145
rect -310 -165 -305 -155
rect -294 -165 -290 -155
rect -310 -175 -290 -165
rect -310 -185 -305 -175
rect -294 -185 -290 -175
rect -310 -195 -290 -185
rect -310 -205 -305 -195
rect -294 -205 -290 -195
rect -310 -210 -290 -205
rect -240 -15 -220 -10
rect -240 -25 -235 -15
rect -224 -25 -220 -15
rect -240 -35 -220 -25
rect -240 -45 -235 -35
rect -224 -45 -220 -35
rect -240 -55 -220 -45
rect -200 -50 -190 -30
rect -170 -32 -160 -30
rect -170 -42 -168 -32
rect -170 -50 -160 -42
rect -240 -65 -235 -55
rect -224 -65 -220 -55
rect -240 -75 -220 -65
rect -120 -66 -100 -60
rect -240 -85 -235 -75
rect -224 -85 -220 -75
rect -240 -95 -220 -85
rect -240 -105 -235 -95
rect -224 -105 -220 -95
rect -240 -115 -220 -105
rect -240 -125 -235 -115
rect -224 -125 -220 -115
rect -240 -135 -220 -125
rect -240 -145 -235 -135
rect -224 -145 -220 -135
rect -240 -155 -220 -145
rect -240 -165 -235 -155
rect -224 -165 -220 -155
rect -120 -155 -115 -66
rect -104 -155 -100 -66
rect -120 -160 -100 -155
rect -50 -66 -30 -60
rect -50 -155 -45 -66
rect -34 -155 -30 -66
rect -50 -160 -30 -155
rect 30 -65 50 -60
rect 30 -155 34 -65
rect 45 -155 50 -65
rect 30 -160 50 -155
rect 100 -65 120 -60
rect 100 -155 105 -65
rect 116 -155 120 -65
rect 100 -160 120 -155
rect -240 -175 -220 -165
rect -240 -185 -235 -175
rect -224 -185 -220 -175
rect -240 -195 -220 -185
rect -240 -205 -235 -195
rect -224 -205 -220 -195
rect -240 -210 -220 -205
<< pdiffusion >>
rect -120 99 -100 110
rect -120 89 -115 99
rect -104 89 -100 99
rect -120 79 -100 89
rect -120 69 -115 79
rect -104 69 -100 79
rect -120 59 -100 69
rect -120 49 -115 59
rect -104 49 -100 59
rect -120 39 -100 49
rect -120 29 -115 39
rect -104 29 -100 39
rect -120 20 -100 29
rect -120 10 -115 20
rect -104 10 -100 20
rect -50 104 -30 110
rect -50 15 -45 104
rect -34 15 -30 104
rect -50 10 -30 15
rect 30 105 50 110
rect 30 15 34 105
rect 45 15 50 105
rect 30 10 50 15
rect 100 100 120 110
rect 100 90 105 100
rect 116 90 120 100
rect 100 80 120 90
rect 100 70 105 80
rect 116 70 120 80
rect 100 60 120 70
rect 100 50 105 60
rect 116 50 120 60
rect 100 40 120 50
rect 100 30 105 40
rect 116 30 120 40
rect 100 20 120 30
rect 100 10 105 20
rect 116 10 120 20
rect 180 98 200 110
rect 180 88 185 98
rect 196 88 200 98
rect 180 79 200 88
rect 180 69 185 79
rect 196 69 200 79
rect 180 59 200 69
rect 180 49 185 59
rect 196 49 200 59
rect 180 40 200 49
rect 180 30 185 40
rect 196 30 200 40
rect 180 20 200 30
rect 180 10 185 20
rect 196 10 200 20
rect 250 105 270 110
rect 250 15 255 105
rect 266 15 270 105
rect 250 10 270 15
<< ndcontact >>
rect -168 -42 -160 -32
rect -115 -155 -104 -66
rect -45 -155 -34 -66
rect 34 -155 45 -65
rect 105 -155 116 -65
<< pdcontact >>
rect -115 89 -104 99
rect -115 69 -104 79
rect -115 49 -104 59
rect -115 29 -104 39
rect -115 10 -104 20
rect -45 15 -34 104
rect 34 15 45 105
rect 105 90 116 100
rect 105 70 116 80
rect 105 50 116 60
rect 105 30 116 40
rect 105 10 116 20
rect 185 88 196 98
rect 185 69 196 79
rect 185 49 196 59
rect 185 30 196 40
rect 185 10 196 20
rect 255 15 266 105
<< psubstratepcontact >>
rect -305 -25 -294 -15
rect -305 -45 -294 -35
rect -305 -65 -294 -55
rect -305 -85 -294 -75
rect -305 -105 -294 -95
rect -305 -125 -294 -115
rect -305 -145 -294 -135
rect -305 -165 -294 -155
rect -305 -185 -294 -175
rect -305 -205 -294 -195
rect -235 -25 -224 -15
rect -235 -45 -224 -35
rect -235 -65 -224 -55
rect -199 -71 -192 -64
rect -186 -71 -179 -64
rect -172 -71 -165 -64
rect -235 -85 -224 -75
rect -235 -105 -224 -95
rect -235 -125 -224 -115
rect -235 -145 -224 -135
rect -235 -165 -224 -155
rect -235 -185 -224 -175
rect -235 -205 -224 -195
rect -240 -245 -229 -234
rect -218 -245 -207 -234
rect -196 -245 -185 -234
<< nsubstratencontact >>
rect -135 119 -128 126
rect -121 119 -114 126
rect -107 119 -100 126
rect -93 119 -86 126
rect -79 119 -72 126
rect -65 119 -58 126
rect -51 119 -44 126
rect -37 119 -30 126
rect -23 119 -16 126
rect 15 119 22 126
rect 29 119 36 126
rect 43 119 50 126
rect 57 119 64 126
rect 71 119 78 126
rect 85 119 92 126
rect 99 119 106 126
rect 113 119 120 126
rect 127 119 134 126
rect 167 119 174 126
rect 181 119 188 126
rect 195 119 202 126
rect 209 119 216 126
rect 223 119 230 126
rect 237 119 244 126
rect 251 119 258 126
rect 265 119 272 126
<< polysilicon >>
rect -100 110 -50 115
rect 50 110 100 115
rect 200 110 250 115
rect -100 8 -50 10
rect 50 8 100 10
rect 200 8 250 10
rect -290 -10 -240 0
rect -190 -29 -185 -25
rect -174 -29 -170 -25
rect -190 -30 -170 -29
rect -190 -55 -170 -50
rect -100 -60 -50 -57
rect 50 -60 100 -48
rect -100 -161 -50 -160
rect 50 -161 100 -160
rect -290 -212 -240 -210
rect -290 -220 -287 -212
rect -241 -220 -240 -212
<< polycontact >>
rect -100 4 -50 8
rect 50 4 100 8
rect 200 1 250 8
rect -185 -29 -174 -25
rect -100 -57 -50 -48
rect -100 -165 -50 -161
rect 50 -165 100 -161
rect -287 -220 -241 -212
<< metal1 >>
rect -128 119 -121 126
rect -114 119 -107 126
rect -100 119 -93 126
rect -86 119 -79 126
rect -72 119 -65 126
rect -58 119 -51 126
rect -44 119 -37 126
rect -30 119 -23 126
rect -16 119 15 126
rect 22 119 29 126
rect 36 119 43 126
rect 50 119 57 126
rect 64 119 71 126
rect 78 119 85 126
rect 92 119 99 126
rect 106 119 113 126
rect 120 119 127 126
rect 134 119 167 126
rect 174 119 181 126
rect 188 119 195 126
rect 202 119 209 126
rect 216 119 223 126
rect 230 119 237 126
rect 244 119 251 126
rect 258 119 265 126
rect 272 119 287 126
rect -115 99 -104 119
rect -115 79 -104 89
rect -115 59 -104 69
rect -115 39 -104 49
rect -305 17 -294 26
rect -115 20 -104 29
rect -305 6 -174 17
rect -305 -15 -294 6
rect -305 -35 -294 -25
rect -305 -55 -294 -45
rect -305 -75 -294 -65
rect -305 -95 -294 -85
rect -305 -115 -294 -105
rect -305 -135 -294 -125
rect -305 -155 -294 -145
rect -305 -175 -294 -165
rect -305 -195 -294 -185
rect -235 -15 -224 -14
rect -235 -35 -224 -25
rect -185 -25 -174 6
rect -235 -55 -224 -45
rect -45 -47 -34 15
rect -100 -48 -34 -47
rect -50 -57 -34 -48
rect -235 -75 -224 -65
rect -45 -66 -34 -57
rect -235 -95 -224 -85
rect -235 -115 -224 -105
rect -235 -135 -224 -125
rect -235 -155 -224 -145
rect -235 -175 -224 -165
rect -235 -195 -224 -185
rect 34 -31 45 15
rect 105 100 116 119
rect 105 80 116 90
rect 105 60 116 70
rect 105 40 116 50
rect 105 20 116 30
rect 185 98 196 119
rect 185 79 196 88
rect 185 59 196 69
rect 185 40 196 49
rect 185 20 196 30
rect 255 105 266 107
rect 214 -31 234 1
rect 255 -6 266 15
rect 34 -38 234 -31
rect 34 -65 45 -38
rect -115 -190 -104 -155
rect 105 -190 116 -155
rect -235 -234 -224 -205
rect -229 -245 -218 -234
rect -207 -245 -196 -234
<< metal2 >>
rect -104 4 100 8
rect -86 -32 -72 4
rect -4 -20 3 4
rect -4 -27 45 -20
rect -199 -64 -191 -34
rect -168 -42 -72 -32
rect -199 -71 -165 -64
rect -100 -165 100 -161
rect -47 -210 -33 -165
rect -287 -220 -33 -210
<< labels >>
rlabel metal1 68 122 68 122 1 Vdd
rlabel metal1 -202 -239 -202 -239 1 gnd
rlabel metal1 -301 12 -301 12 1 d
rlabel metal1 -110 -178 -110 -178 1 a
rlabel metal1 110 -176 110 -176 1 b
rlabel metal1 261 2 261 2 1 vref
<< end >>
