* SPICE3 file created from res2.ext - technology: scmos

.option scale=0.1u

xR0 a 0 b 0 nwellResistor w=12 l=103

.subckt nwellResistor d g s b W=1 L=1 Rsquare = 929
R       d s 'L*Rsquare/W'
Rg      d g 0
Rb      b 0 0
.ends


v a b dc 1.8

.tran 1n 5u
.control
 run
 plot v(a)
.endc
.end
