* SPICE3 file created from bgr1.ext - technology: scmos

.option scale=0.1u

Q1000 0 0 N006 PNP
Q1001 0 0 vctat PNP
Q1002 0 0 N007 PNP
Q1003 0 0 N007 PNP
Q1004 0 0 N007 PNP
Q1005 0 0 N007 PNP
Q1006 0 0 N007 PNP
Q1007 0 0 N007 PNP
Q1008 0 0 N007 PNP
Q1009 0 0 N007 PNP
M1010 N001 N002 N002 N001 pfet w=100 l=50
+  ad=1923.08 pd=230.769 as=1785.71 ps=214.286
Q1011 0 N001 N001 PNP
M1012 0 N003 N004 0 nfet w=200 l=50
+  ad=19400 pd=3936.36 as=3909.43 ps=460.377
M1013 N003 N003 N006 0 nfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240
M1014 N005 N003 N002 0 nfet w=100 l=50
+  ad=1892.86 pd=253.571 as=1916.67 ps=258.333
M1015 N002 N004 0 0 nfet w=20 l=20
+  ad=383.333 pd=51.6667 as=1940 ps=393.636
R0 N005 N007 nwellResistor w=12 l=103
Q1016 0 N001 vref PNP
M1017 N001 N002 vref N001 pfet w=100 l=50
+  ad=1923.08 pd=230.769 as=1785.71 ps=214.286
R1 N001 N004 nwellResistor w=12 l=15428
R2 vref vctat nwellResistor w=12 l=1275
Q1018 0 N001 N002 PNP
M1019 N003 N002 N001 N001 pfet w=100 l=50
+  ad=2000 pd=240 as=1923.08 ps=230.769
C0 N002 N001 7.36fF
C1 N004 0 2.57fF
C2 N003 0 8.80fF
C3 N001 0 61.60fF
C4 N007 0 12.42fF
