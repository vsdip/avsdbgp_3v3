Post Layout Startup Voltage variation

.option scale=0.1u

M1000 N002 N002 N001 N001 pfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240

M1001 N004 N003 0 0 nfet w=200 l=50
+  ad=6000 pd=1300 as=3909.43 ps=460.377

M1002 N006 N003 N003 0 nfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240

M1003 N002 N003 N005 0 nfet w=100 l=50
+  ad=1892.86 pd=253.571 as=1916.67 ps=258.333

M1004 0 N004 N002 0 nfet w=20 l=20
+  ad=383.333 pd=51.6667 as=600 ps=130


M1005 vref N002 N001 N001 pfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240


M1006 N001 N002 N003 N001 pfet w=100 l=50
+  ad=2000 pd=240 as=2000 ps=240


xR0 N005 N007 nwellResistor w=12 l=103
xR1 N001 N004 nwellResistor w=12 l=15428
xR2 vref vctat nwellResistor w=12 l=1275



C0 N001 N002 7.36fF
C1 N004 0 2.57fF
C2 N003 0 8.80fF
C3 N001 0 58.37fF

V1 N001 0 dc pulse 0 3.3 0 50u 50u 1 2
R4 vref 0 100Meg

Q1 0 0 N006 0 2NN2907
Q2 0 0 N007 0 2NN2907 8
Q3 0 0 vctat 0 2NN2907

.MODEL nfet NMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 2.3549E17      VTH0    = 0.3662473
+K1      = 0.5864999      K2      = 1.127266E-3    K3      = 1E-3
+K3B     = 0.0294061      W0      = 1E-7           NLX     = 1.630684E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 1.2064649      DVT1    = 0.4215486      DVT2    = 0.0197749
+U0      = 273.8094484    UA      = -1.40499E-9    UB      = 2.408323E-18
+UC      = 6.504826E-11   VSAT    = 1.355009E5     A0      = 2
+AGS     = 0.4449958      B0      = 1.901075E-7    B1      = 4.99995E-6
+KETA    = -0.0164863     A1      = 3.868769E-4    A2      = 0.4640272
+RDSW    = 123.3376355    PRWG    = 0.5            PRWB    = -0.197728
+WR      = 1              WINT    = 0              LINT    = 1.690044E-8
+DWG     = -4.728719E-9
+DWB     = -2.452411E-9   VOFF    = -0.0948017     NFACTOR = 2.1860065
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 2.230928E-3    ETAB    = 6.028975E-5
+DSUB    = 0.0145467      PCLM    = 1.3822069      PDIBLC1 = 0.1762787
+PDIBLC2 = 1.66653E-3     PDIBLCB = -0.1           DROUT   = 0.7694691
+PSCBE1  = 8.91287E9      PSCBE2  = 7.349607E-9    PVAG    = 1.685917E-3
+DELTA   = 0.01           RSH     = 6.7            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 8.23E-10       CGSO    = 8.23E-10       CGBO    = 1E-12
+CJ      = 9.466429E-4    PB      = 0.8            MJ      = 0.3820266
+CJSW    = 2.608154E-10   PBSW    = 0.8            MJSW    = 0.102322
+CJSWG   = 3.3E-10        PBSWG   = 0.8            MJSWG   = 0.102322
+CF      = 0              PVTH0   = -2.199373E-3   PRDSW   = -0.9368961
+PK2     = 1.593254E-3    WKETA   = -2.880976E-3   LKETA   = 7.165078E-3
+PU0     = 6.777519       PUA     = 5.505418E-12   PUB     = 8.84133E-25
+PVSAT   = 2.006286E3     PETA0   = 1.003159E-4    PKETA   = -6.759277E-3
+NOIMOD=2.0E+00		NOIA=1.3182567385564E+19
+NOIB=144543.977074592 NOIC=-1.24515784572817E-12	EF=0.92 EM=41000000 )


.MODEL pfet PMOS (                                LEVEL   = 49
+VERSION = 3.1            TNOM    = 27             TOX     = 4.1E-9
+XJ      = 1E-7           NCH     = 4.1589E17      VTH0    = -0.3906012
+K1      = 0.5341312      K2      = 0.0395326      K3      = 0
+K3B     = 7.4916211      W0      = 1E-6           NLX     = 1.194072E-7
+DVT0W   = 0              DVT1W   = 0              DVT2W   = 0
+DVT0    = 0.5060555      DVT1    = 0.2423835      DVT2    = 0.1
+U0      = 115.6894042    UA      = 1.573746E-9    UB      = 1.874308E-21
+UC      = -1E-10         VSAT    = 1.130982E5     A0      = 1.9976555
+AGS     = 0.4186945      B0      = 1.949178E-7    B1      = 6.422908E-7
+KETA    = 0.0166345      A1      = 0.4749146      A2      = 0.300003
+RDSW    = 198.321294     PRWG    = 0.5            PRWB    = -0.4986647
+WR      = 1              WINT    = 0              LINT    = 2.94454E-8
+DWG     = -2.798724E-8
+DWB     = -4.83797E-10   VOFF    = -0.095236      NFACTOR = 2
+CIT     = 0              CDSC    = 2.4E-4         CDSCD   = 0
+CDSCB   = 0              ETA0    = 1.035504E-3    ETAB    = -4.358398E-4
+DSUB    = 1.816555E-3    PCLM    = 1.3299898      PDIBLC1 = 1.766563E-3
+PDIBLC2 = 7.728395E-7    PDIBLCB = -1E-3          DROUT   = 1.011891E-3
+PSCBE1  = 4.872184E10    PSCBE2  = 5E-10          PVAG    = 0.0209921
+DELTA   = 0.01           RSH     = 7.7            MOBMOD  = 1
+PRT     = 0              UTE     = -1.5           KT1     = -0.11
+KT1L    = 0              KT2     = 0.022          UA1     = 4.31E-9
+UB1     = -7.61E-18      UC1     = -5.6E-11       AT      = 3.3E4
+WL      = 0              WLN     = 1              WW      = 0
+WWN     = 1              WWL     = 0              LL      = 0
+LLN     = 1              LW      = 0              LWN     = 1
+LWL     = 0              CAPMOD  = 2              XPART   = 0.5
+CGDO    = 6.35E-10       CGSO    = 6.35E-10       CGBO    = 1E-12
+CJ      = 1.144521E-3    PB      = 0.8468686      MJ      = 0.4099522
+CJSW    = 2.490749E-10   PBSW    = 0.8769118      MJSW    = 0.3478565
+CJSWG   = 4.22E-10       PBSWG   = 0.8769118      MJSWG   = 0.3478565
+CF      = 0              PVTH0   = 2.302018E-3    PRDSW   = 9.0575312
+PK2     = 1.821914E-3    WKETA   = 0.0222457      LKETA   = -1.495872E-3
+PU0     = -1.5580645     PUA     = -6.36889E-11   PUB     = 1E-21
+PVSAT   = 49.8420442     PETA0   = 2.827793E-5    PKETA   = -2.536564E-3 
+ NOIMOD=2.0E+00		NOIA=3.57456993317604E+18		NOIB=2500
+ NOIC=2.61260020285845E-11	EF=1.1388				EM=41000000 )


.model 2NN2907 PNP(IS=1E-14 VAF=120
+   BF=250 IKF=0.3 XTB=1.5 BR=3
+   CJC=8E-12 CJE=30E-12 TR=100E-9 TF=400E-12
+   ITF=1 VTF=2 XTF=3 RB=10 RC=.3 RE=.2 )


.subckt nwellResistor d s W=1 L=1 Rsquare = 929
R       d s 'L*Rsquare/W'

.ends

.tran 0.1u 500u


.control
 run
 plot v(N001) v(vref) 
.endc
.end
