magic
tech scmos
timestamp 1594647612
<< nwell >>
rect -140 -20 -10 145
rect 40 -20 170 145
rect 220 -20 350 145
<< ntransistor >>
rect -181 -74 -161 -54
rect -280 -304 -230 -104
rect -100 -204 -50 -104
rect 80 -204 130 -104
<< ptransistor >>
rect -100 10 -50 110
rect 80 10 130 110
rect 260 10 310 110
<< ndiffusion >>
rect -196 -59 -181 -54
rect -196 -69 -194 -59
rect -184 -69 -181 -59
rect -196 -74 -181 -69
rect -161 -59 -146 -54
rect -161 -69 -158 -59
rect -148 -69 -146 -59
rect -161 -74 -146 -69
rect -300 -119 -280 -104
rect -300 -129 -295 -119
rect -285 -129 -280 -119
rect -300 -139 -280 -129
rect -300 -149 -295 -139
rect -285 -149 -280 -139
rect -300 -159 -280 -149
rect -300 -169 -295 -159
rect -285 -169 -280 -159
rect -300 -179 -280 -169
rect -300 -189 -295 -179
rect -285 -189 -280 -179
rect -300 -199 -280 -189
rect -300 -209 -295 -199
rect -285 -209 -280 -199
rect -300 -219 -280 -209
rect -300 -229 -295 -219
rect -285 -229 -280 -219
rect -300 -239 -280 -229
rect -300 -249 -295 -239
rect -285 -249 -280 -239
rect -300 -269 -280 -249
rect -300 -279 -295 -269
rect -285 -279 -280 -269
rect -300 -284 -280 -279
rect -300 -294 -295 -284
rect -285 -294 -280 -284
rect -300 -304 -280 -294
rect -230 -119 -210 -104
rect -230 -129 -225 -119
rect -215 -129 -210 -119
rect -230 -139 -210 -129
rect -230 -149 -225 -139
rect -215 -149 -210 -139
rect -230 -159 -210 -149
rect -230 -169 -225 -159
rect -215 -169 -210 -159
rect -230 -179 -210 -169
rect -230 -189 -225 -179
rect -215 -189 -210 -179
rect -230 -199 -210 -189
rect -230 -209 -225 -199
rect -215 -209 -210 -199
rect -120 -123 -100 -104
rect -120 -133 -115 -123
rect -105 -133 -100 -123
rect -120 -143 -100 -133
rect -120 -153 -115 -143
rect -105 -153 -100 -143
rect -120 -163 -100 -153
rect -120 -173 -115 -163
rect -105 -173 -100 -163
rect -120 -183 -100 -173
rect -120 -193 -115 -183
rect -105 -193 -100 -183
rect -120 -204 -100 -193
rect -50 -124 -30 -104
rect -50 -134 -45 -124
rect -35 -134 -30 -124
rect -50 -144 -30 -134
rect -50 -154 -45 -144
rect -35 -154 -30 -144
rect -50 -164 -30 -154
rect -50 -174 -45 -164
rect -35 -174 -30 -164
rect -50 -184 -30 -174
rect -50 -194 -45 -184
rect -35 -194 -30 -184
rect -50 -204 -30 -194
rect 60 -122 80 -104
rect 60 -132 65 -122
rect 75 -132 80 -122
rect 60 -142 80 -132
rect 60 -152 65 -142
rect 75 -152 80 -142
rect 60 -162 80 -152
rect 60 -172 65 -162
rect 75 -172 80 -162
rect 60 -182 80 -172
rect 60 -192 65 -182
rect 75 -192 80 -182
rect 60 -204 80 -192
rect 130 -109 150 -104
rect 130 -119 135 -109
rect 145 -119 150 -109
rect 130 -129 150 -119
rect 130 -139 135 -129
rect 145 -139 150 -129
rect 130 -149 150 -139
rect 130 -159 135 -149
rect 145 -159 150 -149
rect 130 -169 150 -159
rect 130 -179 135 -169
rect 145 -179 150 -169
rect 130 -189 150 -179
rect 130 -199 135 -189
rect 145 -199 150 -189
rect 130 -204 150 -199
rect -230 -219 -210 -209
rect -230 -229 -225 -219
rect -215 -229 -210 -219
rect -230 -239 -210 -229
rect -230 -249 -225 -239
rect -215 -249 -210 -239
rect -230 -264 -210 -249
rect -230 -274 -225 -264
rect -215 -274 -210 -264
rect -230 -284 -210 -274
rect -230 -294 -225 -284
rect -215 -294 -210 -284
rect -230 -304 -210 -294
<< pdiffusion >>
rect -120 108 -100 110
rect -120 98 -115 108
rect -105 98 -100 108
rect -120 88 -100 98
rect -120 78 -115 88
rect -105 78 -100 88
rect -120 68 -100 78
rect -120 58 -115 68
rect -105 58 -100 68
rect -120 48 -100 58
rect -120 38 -115 48
rect -105 38 -100 48
rect -120 28 -100 38
rect -120 18 -115 28
rect -105 18 -100 28
rect -120 10 -100 18
rect -50 105 -30 110
rect -50 95 -45 105
rect -35 95 -30 105
rect -50 85 -30 95
rect -50 75 -45 85
rect -35 75 -30 85
rect -50 65 -30 75
rect -50 55 -45 65
rect -35 55 -30 65
rect -50 45 -30 55
rect -50 35 -45 45
rect -35 35 -30 45
rect -50 25 -30 35
rect -50 15 -45 25
rect -35 15 -30 25
rect -50 10 -30 15
rect 60 105 80 110
rect 60 95 65 105
rect 75 95 80 105
rect 60 85 80 95
rect 60 75 65 85
rect 75 75 80 85
rect 60 65 80 75
rect 60 55 65 65
rect 75 55 80 65
rect 60 45 80 55
rect 60 35 65 45
rect 75 35 80 45
rect 60 25 80 35
rect 60 15 65 25
rect 75 15 80 25
rect 60 10 80 15
rect 130 108 150 110
rect 130 98 135 108
rect 145 98 150 108
rect 130 88 150 98
rect 130 78 135 88
rect 145 78 150 88
rect 130 68 150 78
rect 130 58 135 68
rect 145 58 150 68
rect 130 48 150 58
rect 130 38 135 48
rect 145 38 150 48
rect 130 28 150 38
rect 130 18 135 28
rect 145 18 150 28
rect 130 10 150 18
rect 240 104 260 110
rect 240 94 245 104
rect 255 94 260 104
rect 240 84 260 94
rect 240 74 245 84
rect 255 74 260 84
rect 240 64 260 74
rect 240 54 245 64
rect 255 54 260 64
rect 240 44 260 54
rect 240 34 245 44
rect 255 34 260 44
rect 240 25 260 34
rect 240 15 245 25
rect 255 15 260 25
rect 240 10 260 15
rect 310 108 330 110
rect 310 98 317 108
rect 327 98 330 108
rect 310 88 330 98
rect 310 78 317 88
rect 327 78 330 88
rect 310 68 330 78
rect 310 58 317 68
rect 327 58 330 68
rect 310 48 330 58
rect 310 38 317 48
rect 327 38 330 48
rect 310 28 330 38
rect 310 18 317 28
rect 327 18 330 28
rect 310 10 330 18
<< ndcontact >>
rect -194 -69 -184 -59
rect -158 -69 -148 -59
rect -295 -129 -285 -119
rect -295 -149 -285 -139
rect -295 -169 -285 -159
rect -295 -189 -285 -179
rect -295 -209 -285 -199
rect -295 -229 -285 -219
rect -295 -249 -285 -239
rect -295 -279 -285 -269
rect -295 -294 -285 -284
rect -225 -129 -215 -119
rect -225 -149 -215 -139
rect -225 -169 -215 -159
rect -225 -189 -215 -179
rect -225 -209 -215 -199
rect -115 -133 -105 -123
rect -115 -153 -105 -143
rect -115 -173 -105 -163
rect -115 -193 -105 -183
rect -45 -134 -35 -124
rect -45 -154 -35 -144
rect -45 -174 -35 -164
rect -45 -194 -35 -184
rect 65 -132 75 -122
rect 65 -152 75 -142
rect 65 -172 75 -162
rect 65 -192 75 -182
rect 135 -119 145 -109
rect 135 -139 145 -129
rect 135 -159 145 -149
rect 135 -179 145 -169
rect 135 -199 145 -189
rect -225 -229 -215 -219
rect -225 -249 -215 -239
rect -225 -274 -215 -264
rect -225 -294 -215 -284
<< pdcontact >>
rect -115 98 -105 108
rect -115 78 -105 88
rect -115 58 -105 68
rect -115 38 -105 48
rect -115 18 -105 28
rect -45 95 -35 105
rect -45 75 -35 85
rect -45 55 -35 65
rect -45 35 -35 45
rect -45 15 -35 25
rect 65 95 75 105
rect 65 75 75 85
rect 65 55 75 65
rect 65 35 75 45
rect 65 15 75 25
rect 135 98 145 108
rect 135 78 145 88
rect 135 58 145 68
rect 135 38 145 48
rect 135 18 145 28
rect 245 94 255 104
rect 245 74 255 84
rect 245 54 255 64
rect 245 34 255 44
rect 245 15 255 25
rect 317 98 327 108
rect 317 78 327 88
rect 317 58 327 68
rect 317 38 327 48
rect 317 18 327 28
<< psubstratepcontact >>
rect -987 -428 -977 -418
rect -937 -428 -927 -418
rect -886 -428 -876 -418
rect -836 -428 -826 -418
rect -786 -428 -776 -418
rect -736 -428 -726 -418
rect -684 -428 -674 -418
rect -634 -428 -624 -418
rect -584 -428 -574 -418
rect -534 -428 -524 -418
rect -484 -428 -474 -418
rect -424 -428 -414 -418
rect -374 -428 -364 -418
rect -324 -428 -314 -418
rect -274 -428 -264 -418
rect -224 -428 -214 -418
rect -174 -428 -164 -418
rect -124 -428 -114 -418
rect -74 -428 -64 -418
rect -24 -428 -14 -418
rect 26 -428 36 -418
rect 76 -428 86 -418
rect 126 -428 136 -418
rect 176 -428 186 -418
rect 226 -428 236 -418
rect 276 -428 286 -418
rect 326 -428 336 -418
rect 376 -428 386 -418
rect 426 -428 436 -418
rect 476 -428 486 -418
rect 526 -428 536 -418
rect 576 -428 586 -418
rect 626 -428 636 -418
rect 676 -428 686 -418
rect 726 -428 736 -418
rect 786 -428 796 -418
rect 836 -428 846 -418
<< nsubstratencontact >>
rect -104 131 -93 141
rect -65 131 -54 141
rect -34 131 -23 141
rect 52 131 63 141
rect 77 131 88 141
rect 106 131 117 141
rect 135 131 146 141
rect 236 131 247 141
rect 269 131 280 141
rect 299 131 310 141
rect -970 119 -958 131
rect 245 -65 257 -53
rect -410 -265 -398 -253
rect -974 -284 -964 -274
rect -944 -284 -934 -274
rect -914 -284 -904 -274
rect -884 -284 -874 -274
rect -854 -284 -844 -274
rect -824 -284 -814 -274
rect -794 -284 -784 -274
rect -764 -284 -754 -274
rect -734 -284 -724 -274
rect -704 -284 -694 -274
rect -674 -284 -664 -274
rect -644 -284 -634 -274
rect -614 -284 -604 -274
rect -584 -284 -574 -274
rect -554 -284 -544 -274
rect -524 -284 -514 -274
rect -494 -284 -484 -274
rect -464 -284 -454 -274
rect -434 -284 -424 -274
rect 356 -129 368 -117
rect 289 -149 299 -139
rect 314 -149 324 -139
rect 135 -258 145 -246
rect 248 -258 258 -246
rect 154 -274 164 -264
rect 193 -274 203 -264
<< polysilicon >>
rect -100 123 -50 125
rect -100 113 -95 123
rect -85 113 -72 123
rect -62 113 -50 123
rect -100 110 -50 113
rect 80 123 130 125
rect 80 113 87 123
rect 97 113 108 123
rect 118 113 130 123
rect 80 110 130 113
rect 260 123 310 125
rect 260 113 265 123
rect 275 113 285 123
rect 295 113 310 123
rect 260 110 310 113
rect -100 -5 -50 10
rect 80 -5 130 10
rect 260 -6 310 10
rect -181 -41 -161 -39
rect -181 -51 -176 -41
rect -166 -51 -161 -41
rect -181 -54 -161 -51
rect -181 -89 -161 -74
rect -280 -92 -230 -89
rect -280 -102 -272 -92
rect -262 -102 -250 -92
rect -240 -102 -230 -92
rect -280 -104 -230 -102
rect -100 -92 -50 -89
rect -100 -102 -95 -92
rect -85 -102 -72 -92
rect -62 -102 -50 -92
rect -100 -104 -50 -102
rect 80 -104 130 -89
rect -100 -207 -50 -204
rect -100 -217 -93 -207
rect -83 -217 -67 -207
rect -57 -217 -50 -207
rect -100 -219 -50 -217
rect 80 -207 130 -204
rect 80 -217 86 -207
rect 96 -217 109 -207
rect 119 -217 130 -207
rect 80 -219 130 -217
rect -280 -319 -230 -304
<< polycontact >>
rect -95 113 -85 123
rect -72 113 -62 123
rect 87 113 97 123
rect 108 113 118 123
rect 265 113 275 123
rect 285 113 295 123
rect -176 -51 -166 -41
rect -272 -102 -262 -92
rect -250 -102 -240 -92
rect -95 -102 -85 -92
rect -72 -102 -62 -92
rect -93 -217 -83 -207
rect -67 -217 -57 -207
rect 86 -217 96 -207
rect 109 -217 119 -207
<< metal1 >>
rect -1010 160 865 170
rect -970 131 -958 160
rect -115 141 -105 160
rect -31 141 -20 160
rect -128 131 -104 141
rect -93 131 -65 141
rect -54 131 -34 141
rect -23 131 -20 141
rect 52 141 63 160
rect 135 141 145 160
rect 233 141 244 160
rect 317 141 327 160
rect 63 131 77 141
rect 88 131 106 141
rect 117 131 135 141
rect 146 131 160 141
rect 233 131 236 141
rect 247 131 269 141
rect 280 131 299 141
rect 310 131 341 141
rect -115 108 -105 131
rect -98 113 -95 123
rect -85 113 -72 123
rect -62 113 87 123
rect 97 113 108 123
rect 118 113 127 123
rect 65 105 75 113
rect -115 88 -105 98
rect -115 68 -105 78
rect -115 48 -105 58
rect -115 28 -105 38
rect -115 13 -105 18
rect -45 85 -35 95
rect -45 65 -35 75
rect -45 45 -35 55
rect -45 25 -35 35
rect -295 -51 -176 -41
rect -166 -51 -163 -41
rect -295 -119 -285 -51
rect -194 -59 -184 -58
rect -159 -69 -158 -59
rect -148 -69 -141 -59
rect -194 -74 -184 -69
rect -275 -102 -272 -92
rect -262 -102 -250 -92
rect -240 -102 -95 -92
rect -85 -102 -72 -92
rect -62 -102 -55 -92
rect -295 -139 -285 -129
rect -295 -159 -285 -149
rect -295 -179 -285 -169
rect -295 -199 -285 -189
rect -295 -219 -285 -209
rect -295 -239 -285 -229
rect -295 -253 -285 -249
rect -398 -265 -285 -253
rect -295 -269 -285 -265
rect -998 -284 -974 -274
rect -964 -284 -944 -274
rect -934 -284 -914 -274
rect -904 -284 -884 -274
rect -874 -284 -854 -274
rect -844 -284 -824 -274
rect -814 -284 -794 -274
rect -784 -284 -764 -274
rect -754 -284 -734 -274
rect -724 -284 -704 -274
rect -694 -284 -674 -274
rect -664 -284 -644 -274
rect -634 -284 -614 -274
rect -604 -284 -584 -274
rect -574 -284 -554 -274
rect -544 -284 -524 -274
rect -514 -284 -494 -274
rect -484 -284 -464 -274
rect -454 -284 -434 -274
rect -424 -284 -371 -274
rect -295 -284 -285 -279
rect -997 -418 -987 -284
rect -684 -418 -674 -284
rect -389 -418 -379 -284
rect -295 -299 -285 -294
rect -225 -119 -215 -109
rect -225 -139 -215 -129
rect -225 -159 -215 -149
rect -225 -179 -215 -169
rect -225 -199 -215 -189
rect -225 -219 -215 -209
rect -225 -239 -215 -229
rect -225 -264 -215 -249
rect -115 -123 -105 -109
rect -115 -143 -105 -133
rect -115 -163 -105 -153
rect -115 -183 -105 -173
rect -115 -253 -105 -193
rect -45 -124 -35 15
rect 65 85 75 95
rect 65 65 75 75
rect 65 45 75 55
rect 65 25 75 35
rect 65 3 75 15
rect 135 108 145 131
rect 251 113 265 123
rect 275 113 285 123
rect 295 113 306 123
rect 317 108 327 131
rect 135 88 145 98
rect 135 68 145 78
rect 135 48 145 58
rect 135 28 145 38
rect 135 13 145 18
rect 245 104 255 106
rect 245 84 255 94
rect 245 64 255 74
rect 245 44 255 54
rect 245 25 255 34
rect 245 -53 255 15
rect 317 88 327 98
rect 317 68 327 78
rect 317 48 327 58
rect 317 28 327 38
rect 317 13 327 18
rect 582 59 874 69
rect 582 7 592 59
rect 729 26 760 35
rect 582 -3 642 7
rect 738 -3 748 26
rect 864 7 874 59
rect 840 -3 874 7
rect -45 -144 -35 -134
rect -45 -164 -35 -154
rect -45 -184 -35 -174
rect -45 -207 -35 -194
rect 65 -122 75 -99
rect 582 -99 592 -3
rect 729 -12 760 -3
rect 738 -71 748 -12
rect 729 -80 760 -71
rect 582 -109 642 -99
rect 65 -142 75 -132
rect 65 -162 75 -152
rect 65 -182 75 -172
rect 65 -197 75 -192
rect 135 -129 145 -119
rect 135 -149 145 -139
rect 287 -149 289 -139
rect 299 -149 314 -139
rect 324 -149 339 -139
rect 135 -169 145 -159
rect 135 -189 145 -179
rect -95 -217 -93 -207
rect -83 -217 -67 -207
rect -57 -217 86 -207
rect 96 -217 109 -207
rect 119 -217 126 -207
rect 135 -246 145 -199
rect 137 -274 154 -264
rect 164 -274 193 -264
rect 203 -274 233 -264
rect -225 -284 -215 -274
rect -225 -418 -215 -294
rect -194 -418 -184 -371
rect -105 -418 -96 -340
rect -86 -418 -77 -342
rect 143 -418 153 -274
rect 206 -418 216 -274
rect 248 -336 258 -258
rect 289 -418 299 -149
rect 314 -418 324 -149
rect 356 -159 368 -129
rect 356 -169 381 -159
rect 371 -212 381 -169
rect 582 -205 592 -109
rect 738 -128 748 -80
rect 864 -99 874 -3
rect 840 -109 874 -99
rect 729 -137 760 -128
rect 738 -177 748 -137
rect 728 -186 759 -177
rect 582 -215 642 -205
rect 343 -418 352 -298
rect 381 -418 391 -301
rect 582 -312 592 -215
rect 738 -234 748 -186
rect 864 -205 874 -109
rect 839 -215 874 -205
rect 728 -243 759 -234
rect 738 -284 748 -243
rect 728 -293 759 -284
rect 582 -322 643 -312
rect 582 -356 592 -322
rect 738 -341 748 -293
rect 864 -313 874 -215
rect 843 -323 874 -313
rect 728 -350 759 -341
rect 551 -366 592 -356
rect 738 -418 748 -350
rect -1010 -428 -987 -418
rect -977 -428 -937 -418
rect -927 -428 -886 -418
rect -876 -428 -836 -418
rect -826 -428 -786 -418
rect -776 -428 -736 -418
rect -726 -428 -684 -418
rect -674 -428 -634 -418
rect -624 -428 -584 -418
rect -574 -428 -534 -418
rect -524 -428 -484 -418
rect -474 -428 -424 -418
rect -414 -428 -374 -418
rect -364 -428 -324 -418
rect -314 -428 -274 -418
rect -264 -428 -224 -418
rect -214 -428 -174 -418
rect -164 -428 -124 -418
rect -114 -428 -74 -418
rect -64 -428 -24 -418
rect -14 -428 26 -418
rect 36 -428 76 -418
rect 86 -428 126 -418
rect 136 -428 176 -418
rect 186 -428 226 -418
rect 236 -428 276 -418
rect 286 -428 326 -418
rect 336 -428 376 -418
rect 386 -428 426 -418
rect 436 -428 476 -418
rect 486 -428 526 -418
rect 536 -428 576 -418
rect 586 -428 626 -418
rect 636 -428 676 -418
rect 686 -428 726 -418
rect 736 -428 786 -418
rect 796 -428 836 -418
<< m2contact >>
rect -141 -69 -131 -59
rect -194 -85 -184 -74
rect 241 113 251 123
rect 65 -7 75 3
rect 65 -99 75 -89
rect -194 -371 -184 -361
rect 248 -346 258 -336
rect 541 -366 551 -356
<< metal2 >>
rect 201 113 241 123
rect 65 -59 75 -7
rect -131 -60 75 -59
rect 201 -60 211 113
rect -131 -69 211 -60
rect -194 -361 -184 -85
rect 65 -89 75 -69
rect 248 -356 258 -346
rect 248 -366 541 -356
<< rnwell >>
rect -958 119 -371 131
rect -383 115 -371 119
rect -999 103 -371 115
rect -999 99 -987 103
rect -999 87 -371 99
rect -383 83 -371 87
rect -999 71 -371 83
rect -999 67 -987 71
rect -999 55 -371 67
rect -383 51 -371 55
rect -999 39 -371 51
rect -999 35 -987 39
rect -999 23 -371 35
rect -383 19 -371 23
rect -999 7 -371 19
rect -999 3 -987 7
rect -999 -9 -371 3
rect -383 -13 -371 -9
rect -999 -25 -371 -13
rect -999 -29 -987 -25
rect -999 -41 -371 -29
rect -383 -45 -371 -41
rect -999 -57 -371 -45
rect -999 -61 -987 -57
rect -999 -73 -371 -61
rect -383 -77 -371 -73
rect -999 -89 -371 -77
rect 257 -65 523 -53
rect 511 -69 523 -65
rect -999 -93 -987 -89
rect -999 -105 -371 -93
rect -383 -109 -371 -105
rect -999 -121 -371 -109
rect 221 -81 523 -69
rect 221 -85 233 -81
rect 221 -97 523 -85
rect 511 -101 523 -97
rect -999 -125 -987 -121
rect -999 -137 -371 -125
rect -383 -141 -371 -137
rect -999 -153 -371 -141
rect -999 -157 -987 -153
rect -999 -169 -371 -157
rect -383 -173 -371 -169
rect -999 -185 -371 -173
rect -999 -189 -987 -185
rect -999 -201 -371 -189
rect -383 -205 -371 -201
rect -999 -217 -371 -205
rect -999 -221 -987 -217
rect -999 -233 -371 -221
rect -383 -237 -371 -233
rect -999 -249 -371 -237
rect -999 -253 -987 -249
rect -999 -265 -410 -253
rect 221 -113 523 -101
rect 221 -117 233 -113
rect 221 -129 356 -117
rect 145 -258 248 -246
<< pseudo_nwr >>
rect -1017 131 -353 145
rect -1017 119 -970 131
rect -1017 115 -383 119
rect -1017 87 -999 115
rect -371 103 -353 131
rect -987 99 -353 103
rect -1017 83 -383 87
rect -1017 55 -999 83
rect -371 71 -353 99
rect -987 67 -353 71
rect -1017 51 -383 55
rect -1017 23 -999 51
rect -371 39 -353 67
rect -987 35 -353 39
rect -1017 19 -383 23
rect -1017 -9 -999 19
rect -371 7 -353 35
rect -987 3 -353 7
rect -1017 -13 -383 -9
rect -1017 -41 -999 -13
rect -371 -25 -353 3
rect -987 -29 -353 -25
rect -1017 -45 -383 -41
rect -1017 -73 -999 -45
rect -371 -57 -353 -29
rect 215 -53 529 -42
rect -987 -61 -353 -57
rect -1017 -77 -383 -73
rect -1017 -105 -999 -77
rect -371 -89 -353 -61
rect 215 -65 245 -53
rect 215 -69 511 -65
rect -987 -93 -353 -89
rect -1017 -109 -383 -105
rect -1017 -137 -999 -109
rect -371 -121 -353 -93
rect 215 -97 221 -69
rect 523 -81 529 -53
rect 233 -85 529 -81
rect 215 -101 511 -97
rect -987 -125 -353 -121
rect -1017 -141 -383 -137
rect -1017 -169 -999 -141
rect -371 -153 -353 -125
rect -987 -157 -353 -153
rect -1017 -173 -383 -169
rect -1017 -201 -999 -173
rect -371 -185 -353 -157
rect -987 -189 -353 -185
rect -1017 -205 -383 -201
rect -1017 -233 -999 -205
rect -371 -217 -353 -189
rect -987 -221 -353 -217
rect -1017 -237 -383 -233
rect -1017 -265 -999 -237
rect -371 -249 -353 -221
rect -987 -253 -353 -249
rect -398 -265 -353 -253
rect -1017 -274 -353 -265
rect -1017 -284 -974 -274
rect -964 -284 -944 -274
rect -934 -284 -914 -274
rect -904 -284 -884 -274
rect -874 -284 -854 -274
rect -844 -284 -824 -274
rect -814 -284 -794 -274
rect -784 -284 -764 -274
rect -754 -284 -734 -274
rect -724 -284 -704 -274
rect -694 -284 -674 -274
rect -664 -284 -644 -274
rect -634 -284 -614 -274
rect -604 -284 -584 -274
rect -574 -284 -554 -274
rect -544 -284 -524 -274
rect -514 -284 -494 -274
rect -484 -284 -464 -274
rect -454 -284 -434 -274
rect -424 -284 -353 -274
rect -1017 -285 -353 -284
rect 215 -129 221 -101
rect 523 -113 529 -85
rect 233 -117 529 -113
rect 368 -129 529 -117
rect 215 -139 529 -129
rect 215 -149 289 -139
rect 299 -149 314 -139
rect 324 -149 529 -139
rect 215 -158 529 -149
rect 125 -246 279 -236
rect 125 -258 135 -246
rect 258 -258 279 -246
rect 125 -264 279 -258
rect 125 -274 154 -264
rect 164 -274 193 -264
rect 203 -274 279 -264
rect 125 -278 279 -274
use p  p_0
timestamp 1594489297
transform 1 0 -157 0 1 -331
box 5 -13 89 79
use p  p_1
timestamp 1594489297
transform 1 0 329 0 1 -290
box 5 -13 89 79
use p  p_2
timestamp 1594489297
transform 0 -1 719 1 0 -257
box 5 -13 89 79
use p  p_3
timestamp 1594489297
transform 0 -1 719 1 0 -364
box 5 -13 89 79
use p  p_4
timestamp 1594489297
transform 0 1 767 -1 0 -163
box 5 -13 89 79
use p  p_5
timestamp 1594489297
transform 0 1 767 -1 0 -270
box 5 -13 89 79
use p  p_6
timestamp 1594489297
transform 0 -1 719 1 0 -151
box 5 -13 89 79
use p  p_7
timestamp 1594489297
transform 0 -1 719 1 0 -45
box 5 -13 89 79
use p  p_9
timestamp 1594489297
transform 0 1 767 -1 0 49
box 5 -13 89 79
use p  p_8
timestamp 1594489297
transform 0 1 767 -1 0 -57
box 5 -13 89 79
<< labels >>
rlabel metal1 13 117 13 117 1 N002
rlabel metal1 -41 -47 -41 -47 1 N003
rlabel metal1 -350 -261 -350 -261 1 N004
rlabel metal1 140 -227 140 -227 1 N005
rlabel metal1 -110 -206 -110 -206 1 N006
rlabel metal1 247 -31 247 -31 1 vref
rlabel metal1 364 -157 364 -157 1 vctat
rlabel metal1 -27 -423 -27 -423 1 0
rlabel metal1 -55 164 -55 164 1 N001
rlabel metal1 253 -279 253 -279 1 N007
<< end >>
