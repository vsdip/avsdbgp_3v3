magic
tech scmos
timestamp 1593461626
<< nwell >>
rect -31 -29 31 29
<< pdiffusion >>
rect -20 16 20 18
rect -20 12 -14 16
rect -10 12 -3 16
rect 1 12 9 16
rect 13 12 20 16
rect -20 10 20 12
rect -20 6 -18 10
rect -14 6 -12 10
rect 12 6 14 10
rect 18 6 20 10
rect -20 2 -12 6
rect -20 -2 -18 2
rect -14 -2 -12 2
rect -20 -6 -12 -2
rect -8 2 8 6
rect -8 -2 -2 2
rect 2 -2 8 2
rect -8 -6 8 -2
rect 12 2 20 6
rect 12 -2 14 2
rect 18 -2 20 2
rect 12 -6 20 -2
rect -20 -10 -18 -6
rect -14 -10 -12 -6
rect 12 -10 14 -6
rect 18 -10 20 -6
rect -20 -12 20 -10
rect -20 -16 -14 -12
rect -10 -16 -2 -12
rect 2 -16 10 -12
rect 14 -16 20 -12
rect -20 -18 20 -16
<< pdcontact >>
rect -14 12 -10 16
rect -3 12 1 16
rect 9 12 13 16
rect -18 6 -14 10
rect 14 6 18 10
rect -18 -2 -14 2
rect -2 -2 2 2
rect 14 -2 18 2
rect -18 -10 -14 -6
rect 14 -10 18 -6
rect -14 -16 -10 -12
rect -2 -16 2 -12
rect 10 -16 14 -12
<< psubstratepcontact >>
rect -32 32 -22 37
rect 0 32 10 37
rect 25 32 35 37
rect -40 2 -34 17
rect 34 4 40 19
rect -40 -25 -34 -10
rect 34 -26 40 -11
rect -30 -37 -9 -32
rect 6 -37 27 -32
<< nsubstratencontact >>
rect -28 22 -24 26
rect -20 22 -16 26
rect -12 22 -8 26
rect -4 22 0 26
rect 4 22 8 26
rect 12 22 16 26
rect 20 22 24 26
rect -28 14 -24 18
rect 24 14 28 18
rect -28 6 -24 10
rect 24 6 28 10
rect -28 -2 -24 2
rect 24 -2 28 2
rect -28 -10 -24 -6
rect 24 -10 28 -6
rect -28 -18 -24 -14
rect 24 -18 28 -14
rect -24 -26 -20 -22
rect -14 -26 -10 -22
rect -6 -26 -2 -22
rect 2 -26 6 -22
rect 10 -26 14 -22
rect 18 -26 22 -22
<< metal1 >>
rect -40 32 -32 37
rect -22 32 0 37
rect 10 32 25 37
rect 35 32 40 37
rect -40 17 -34 32
rect -40 -10 -34 2
rect -40 -32 -34 -25
rect -24 22 -20 26
rect -16 22 -12 26
rect -8 22 -4 26
rect 0 22 4 26
rect 8 22 12 26
rect 16 22 20 26
rect -28 18 -24 22
rect 24 18 28 26
rect -28 10 -24 14
rect -28 2 -24 6
rect -28 -6 -24 -2
rect -28 -14 -24 -10
rect -18 10 -14 16
rect -10 12 -3 16
rect 1 12 9 16
rect 13 12 18 16
rect -18 2 -14 6
rect 14 10 18 12
rect -18 -6 -14 -2
rect -5 2 5 4
rect -5 -2 -2 2
rect 2 -2 5 2
rect -5 -4 5 -2
rect 14 2 18 6
rect -18 -16 -14 -10
rect 14 -6 18 -2
rect -10 -16 -2 -12
rect 2 -16 10 -12
rect 14 -16 18 -10
rect 24 10 28 14
rect 24 2 28 6
rect 24 -6 28 -2
rect 24 -14 28 -10
rect -28 -26 -24 -18
rect 24 -22 28 -18
rect -20 -26 -14 -22
rect -10 -26 -6 -22
rect -2 -26 2 -22
rect 6 -26 10 -22
rect 14 -26 18 -22
rect 22 -26 28 -22
rect 34 19 40 32
rect 34 -11 40 4
rect 34 -32 40 -26
rect -40 -37 -30 -32
rect -9 -37 6 -32
rect 27 -37 40 -32
<< labels >>
rlabel metal1 -4 -3 -4 -3 1 e
rlabel metal1 -16 12 -16 12 1 c
rlabel metal1 -22 24 -22 24 1 b
rlabel metal1 38 21 38 21 7 gnd
<< end >>
