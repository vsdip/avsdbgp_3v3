magic
tech scmos
timestamp 1593889714
<< nsubstratencontact >>
rect -31 7 -25 19
rect 31 7 37 19
<< rnwell >>
rect -25 7 31 19
<< pseudo_nwr >>
rect -37 19 41 23
rect -37 7 -31 19
rect 37 7 41 19
rect -37 -17 41 7
<< labels >>
rlabel nsubstratencontact -29 13 -29 13 1 a
rlabel nsubstratencontact 33 13 33 13 1 b
<< end >>
